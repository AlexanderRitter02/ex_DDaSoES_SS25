module fuse (
    input  logic a,
    input  logic set,
    output logic b
);

  // TODO
endmodule
