module and(
  input logic a, b
  output logic o
)

  assign o = a & b

endmodule
