package fourteen_segment_display;

//typedef logic [14 : 0] display_pins_t;

localparam logic [14 : 0] R = 'b001110001001101;
localparam logic [14 : 0] O = 'b001010100010101;
localparam logic [14 : 0] C = 'b001010100000001;
localparam logic [14 : 0] W = 'b001011001010100;
localparam logic [14 : 0] C_dot = 'b001010100100001;
localparam logic [14 : 0] W_dot = 'b001011001110100;

endpackage